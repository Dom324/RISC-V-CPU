module CPU(
  input keyboard_data, keyboard_clock,
  input CLK_VGA, CLK_CPU,
  output hsync, vsync, VGA_pixel
  );


endmodule
